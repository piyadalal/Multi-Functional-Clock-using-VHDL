library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package ddram_package is
	type ddram_x_y is array (0 to 19, 0 to 3) of character;
end ddram_package;